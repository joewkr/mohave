netcdf test3 {
types:
  compound c1 {
    uint a;
    ubyte b;
  }

  compound compound_t {
    int n;
    float x\ field\ name;
    float y;
  }

  compound compound_with_strings {
    int n;
    string comment;
  }

  byte enum qa_flags {Best\ quality = 0, Good\ quality = 1, Poor\ quality = 2, No\ decision= 127};
  short enum precip_type {None = 999, Rain = 0, Snow = 1};

  double(*) profile;
  compound_t(*) compound_profile;

  opaque(65) binary_blob;
  opaque(1) binary_mb;

dimensions:
  dim1 = 3;
  dim2 = 2;
  dim3 = 1;
variables:
  int scalar_int;
    int64 scalar_int:many_ints = 3, 7, 21;
  compound_t scalar_compound;
  compound_t vector_compound(dim1);
  compound_with_strings vector_compound_ws(dim1);
  binary_blob scalar_opaque;
    binary_mb scalar_opaque:attr = 0X00, 0X02;
    binary_mb scalar_opaque:scalar\ attr = 0X01;
  qa_flags scalar_enum;
    precip_type scalar_enum:attr = None, Rain, Snow;
    precip_type scalar_enum:scalar\ attr = Snow;
  qa_flags vector_enum(dim1);
  profile scalar_vlen;
  profile vector_vlen(dim1);
  compound_profile vector_vlen_compound(dim1);
    compound_profile vector_vlen_compound:attr = {{7, 2.54, -7.99}, {1, 2.2, 3.3}}, {{5.5, 6.6, 7.7}};
    compound_profile vector_vlen_compound:scalar\ attr = {{7, 2.54, -7.99}, {1, 2.2, 3.3}, {5.5, 6.6, 7.7}};
  int vector_int(dim1);
  float vector_float(dim1);
  string just_string;
  string string_vector(dim1);
    string string_vector:long_name = "a vector of strings";
    double string_vector:test_attr = 1.5;
  string string_matrix(dim2, dim1);

// global attributes:
  string :summary = "test NetCDF file", "NetCDF4";
  int :version = 2021;
data:
  scalar_int = 7;
  scalar_compound = { 18, 0.2f, 34.56f};
  vector_compound = { 17, 0.1f, 23.45f}, {-1, 22.44f, 1.0e+20}, {22, 1.0f, 5.7f};
  vector_compound_ws = {1, "hello"}, {-1, "world"}, {177, "long comment"};
  scalar_opaque = 0X0123456789ABCDEF0123456789ABCDEF11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010;
  scalar_enum = Poor\ quality;
  vector_enum = No\ decision, Best\ quality, Good\ quality;
  scalar_vlen = {1,2,3,4,6};
  vector_vlen = {1,2}, {9,100,-777}, {22.33, 77.98, 123.789, 0.554};
  vector_vlen_compound = {{7, 57.98f, 12.34f}, {1, 2.0f, 11.75f}}, {{19, 0.2f, 34.56f}}, {{1, -12.22f, -13.54f}, {2, 65.56f, 123.321f}, {0, 0.1f, 0.2f}};
  vector_int = 3, 4, 5;
  vector_float = 13.4f, 14.5f, 15.6f;
  just_string = "some text";
  string_vector = "one", "two", "three";
  string_matrix = "aa", "bb", "cc", "dd", "ee", "ff";
}
