netcdf empty {}
