netcdf test1 {
dimensions:
  dim1 = 7;
  dim2 = 3;
  dim3 = 21;
  dim4 = UNLIMITED;
variables:
  double dummy_var;
    dummy_var:_Endianness = "little";
  float scalar_var;
    scalar_var:_Endianness = "big";
    scalar_var:long_name = "scalar variable";
    scalar_var:units = "m/s";
  int vector_var(dim1);
    vector_var:_DeflateLevel = 9;
    vector_var:_FillValue = 1;
    vector_var:_Fletcher32 = "true";
  int var_2d(dim1, dim2);
    var_2d:_ChunkSizes = 2, 3;
    var_2d:_Shuffle = "true";
  int var_2d_compressed4(dim1, dim2);
    var_2d_compressed4:_ChunkSizes = 2, 3;
    var_2d_compressed4:_Shuffle = "true";
    var_2d_compressed4:_DeflateLevel = 4;
  int var_2d_compressed0(dim1, dim2);
    var_2d_compressed0:_ChunkSizes = 2, 3;
    var_2d_compressed0:_Shuffle = "true";
    var_2d_compressed0:_DeflateLevel = 0;
  int var_unlim(dim4);
}
